module stream_rx(
    // system signals
    input                   sclk,
    input                   s_rst_n,
    // Stream Rx Interface
    input           [63:0]  s_axis_mm2s_tdata,
    input           [ 7:0]  s_axis_mm2s_tkeep, // tkeep Ӧ��Ҳ�����ݣ���ʹδʹ��
    input                   s_axis_mm2s_tvalid,
    output  wire            s_axis_mm2s_tready,
    input                   s_axis_mm2s_tlast,
    // Main Ctrl Interface
    input           [ 1:0]  data_type,
    input           [ 5:0]  state,
    output  wire            write_finish,
    // Output data and valid signals
    output  reg     [63:0]  stream_rx_data,
    output  reg             stream_feature_vld,
    output  reg             stream_weight_vld,
    output  reg             stream_bias_vld,
    output  reg             stream_leakyrelu_vld
);

//========================================================================\
// =========== Define Parameter and Internal signals =========== 
//========================================================================/
localparam      FEATURE_DATA    = 2'b00;
localparam      WEIGHT_DATA     = 2'b01;
localparam      BIAS_DATA       = 2'b10;
localparam      LEAKYRELU_DATA  = 2'b11;

// �ڲ���ˮ�߼Ĵ���
reg             internal_vld;
reg             internal_tlast;
reg     [63:0]  internal_tdata;
reg     [ 1:0]  internal_data_type; // ����data_type�Է������б仯

//=============================================================================
//**************    Main Code   **************
//=============================================================================

// 1. ������ʱ������������
// ����״̬����(state[1]) ���� �ڲ���ˮ��Ϊ����ʱ( !internal_vld )�����ǲ�׼���ý���������
assign  s_axis_mm2s_tready = state[1] & !internal_vld;

// 2. �����������ݵ��ڲ���ˮ�߼Ĵ���
// �����ֳɹ�ʱ (tvalid & tready)�����������ݴ���Ĵ���
always @(posedge sclk or negedge s_rst_n) begin
    if (s_rst_n == 1'b0) begin
        internal_vld <= 1'b0;
    end else if (s_axis_mm2s_tvalid && s_axis_mm2s_tready) begin
        internal_vld <= 1'b1; // ������Ч
        internal_tdata <= s_axis_mm2s_tdata;
        internal_tlast <= s_axis_mm2s_tlast;
        internal_data_type <= data_type; // �����ݰ���ʼʱ��������
    end else begin
        internal_vld <= 1'b0; // �����������ˮ�߱���Ч
    end
end

// 3. ������������ݲ������
// ����ź������ǼĴ������������ȷ��ʱ��
always @(posedge sclk or negedge s_rst_n) begin
    if (s_rst_n == 1'b0) begin
        stream_rx_data <= 64'b0;
        stream_feature_vld <= 1'b0;
        stream_weight_vld <= 1'b0;
        stream_bias_vld <= 1'b0;
        stream_leakyrelu_vld <= 1'b0;
    end else if (internal_vld) begin // ���ڲ��Ĵ�����Чʱ
        stream_rx_data <= internal_tdata;
        // ���������data_type��������Ӧ��vld�ź�
        stream_feature_vld <= (internal_data_type == FEATURE_DATA) ? 1'b1 : 1'b0;
        stream_weight_vld  <= (internal_data_type == WEIGHT_DATA) ? 1'b1 : 1'b0;
        stream_bias_vld    <= (internal_data_type == BIAS_DATA) ? 1'b1 : 1'b0;
        stream_leakyrelu_vld <= (internal_data_type == LEAKYRELU_DATA) ? 1'b1 : 1'b0;
    end else begin
        stream_rx_data <= 64'b0; // Ĭ��ֵ
        stream_feature_vld <= 1'b0;
        stream_weight_vld <= 1'b0;
        stream_bias_vld <= 1'b0;
        stream_leakyrelu_vld <= 1'b0;
    end
end

// 4. write_finish �ź�
// ���ڲ��Ĵ�����Ч�������һ�����ݰ�ʱ����������ź�
assign write_finish = internal_vld & internal_tlast;


endmodule