module LIF #(
    parameter INPUT_WIDTH       = 8,    
    parameter VOLTAGE_WIDTH     = 16,  
    parameter VOLTAGE_FRAC_BITS = 8, 
    // ��ֵ��Ϊ1.0
    parameter THRESHOLD         = 16'h0100 
)(
    // ϵͳ�ź�
    input                           clk,
    input                           rst_n,
    // �����ź�
    input                           i_valid,        // ����������Ч�ź�
    input      signed [INPUT_WIDTH-1:0]   neuron_in,      // �������ݣ����磺���Ծ������ۼӽ����
    // ����ź�
    output     reg                    spike_out,      // ������� (1 ��ʾ����, 0 ��ʾ������)
    output     reg                    o_valid         // ���������Ч�ź�
);

// �ڲ�Ĥ��λ�Ĵ���������Ϊ�з������Դ���������ѹ
reg   signed [VOLTAGE_WIDTH-1:0]    membrane_potential;

wire  signed [VOLTAGE_WIDTH-1:0]    leaky_potential;
wire  signed [VOLTAGE_WIDTH-1:0]    scaled_input;
wire  signed [VOLTAGE_WIDTH-1:0]    next_membrane_potential;

assign leaky_potential = membrane_potential - (membrane_potential >> 2);
assign scaled_input = {{(VOLTAGE_WIDTH-INPUT_WIDTH){neuron_in[INPUT_WIDTH-1]}}, neuron_in};
assign next_membrane_potential = leaky_potential + scaled_input;

//charge  0.25 0.4375 0.5781 0.6836
// def neuronal_charge_decay_input_reset0(x: torch.Tensor, v: torch.Tensor, tau: float):
// v = v + (x - v) / tau
// return v

// --- �ӳٿ����߼� ---
// ����һ�������ӳٵ�������Ч�źţ�����ͬ�����
reg i_valid_d1;
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        i_valid_d1 <= 1'b0;
        o_valid    <= 1'b0;
    end else begin
        i_valid_d1 <= i_valid;
        o_valid <= i_valid_d1;
    end
end


// --- Ĥ��λ�����߼� ---
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        membrane_potential <= 'd0;
        spike_out          <= 1'b0;
    end else begin
        // Ĭ������£��������Ϊ0
        spike_out <= 1'b0;

        if (i_valid_d1) begin // ��������Ч����һ�Ľ��м���
            // �����һ���ڵ�Ĥ��λ�Ƿ񳬹���ֵ
            if (membrane_potential > THRESHOLD) begin
                // A. ���Ų����� (Fire and Reset)
                spike_out          <= 1'b1;   // ��������
                membrane_potential <= 'd0;     // Ĥ��λ����Ϊ0
            end else begin
                // B. й©������ (Leaky and Integrate)
                membrane_potential <= next_membrane_potential;
            end
        end
    end
end

endmodule